module jkflop(clk, j, k, q);
    input clk, j, k;
    output q;

endmodule
