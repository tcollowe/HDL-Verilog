module tflop(q, clk, t);
    input clk, t;
    output q;

endmodule
