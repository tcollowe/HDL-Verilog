`default_nettype none
`timescale 1ns/1ns

module test_mult4();
    wire a, b, c;

    mult4 uut1(a, b, c);
    initial begin
        
    end



endmodule