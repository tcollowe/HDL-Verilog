module tflop(clk, t, q);
    input clk, t;
    output q;

endmodule
