module priority4 (in, out, valid);
	input wire[3:0] in;
	output reg[1:0] out;
	output wire valid;



	
endmodule