/*
Use the XOR primitive and your D-flip-flop to implement the T flipflop:
*/

module tflop(clk, t, q);
    input clk, t;
    output q;

endmodule
