module func(sel,
            x,
            y,
            z);

    input [3:0] sel;
    input x, y;
    output reg z;

    always @() begin
        
    end


    
endmodule
