/*
Implement the S-R latch using two NAND gate primitives using the same logic table as before (not the one shown in the text, or here).  Note: because the truth table is *different* than it is from the textbook, you will need to do more than just include just two NAND gates.  
*/

module srlatch(e, s, r, q);
    input e, s, r;
    inout q;

endmodule

