module jkflop(q, clk, j, k);
    input clk, j, k;
    output q;

endmodule
