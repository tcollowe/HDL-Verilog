module hello();
    
    initial begin
        $display("Hello World\n");
    end
    
endmodule
