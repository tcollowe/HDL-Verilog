`default_nettype none
module mult (a, b, c);
    input wire[3:0] a;
    input wire[3:0] b;
    output wire[7:0] c;
    
endmodule