module dlatch(clk, d, q);
    input clk, d;
    output q;

endmodule
