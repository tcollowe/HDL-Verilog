module dflop(q, clk, d);
    input clk, d;
    output q;

endmodule
