`default_nettype none
module mult4 (a, b, c);
    input wire[3:0] a;
    input wire[3:0] b;
    output wire[7:0] c;
    
endmodule