module dflop(clk, d, q);
    input clk, d;
    output q;

endmodule
