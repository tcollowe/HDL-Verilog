`default_nettype none
`timescale 1ns/1ns

module test_mult();
    wire a, b, c;

    mult uut1(a, b, c);
    initial begin
        
    end



endmodule