`default_nettype none
`timescale 1ns/1ps

module test();

initial begin
	$display("hello world\n");
end

endmodule
